module control_unit (
    input [31:0]   instr,
    output         write_reg,
    output         mem_write,
    output         bus_write,
);
    
endmodule