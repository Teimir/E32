module E32(
   input clk,
	output led
);

endmodule